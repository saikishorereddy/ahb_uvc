module ahb_slave();
endmodule
