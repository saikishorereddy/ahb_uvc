interface ahb_intf(input logic hclk, hrstn);
endinterface
